module NOT(input logic a, output logic b);

assign b = ~a;

endmodule
 
